package state_type_package is
	TYPE State_type is (S0, S1, S2A, S2B, S3, S4);
end package;